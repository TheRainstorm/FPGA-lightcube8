`include "defines.h"

module frame_buffer (
    input wire clk,
    input wire rst,
    input wire [1: 0] display_mode,
    input wire [3: 0] display_sel,

    input wire [8*64-1: 0] frame_cube_uart_flat,
    input wire frame_valid_uart,
    input wire [8*64-1: 0] frame_cube_default_flat,
    input wire frame_valid_default,

    output reg [31: 0] frame_cnt,
    output reg [8*64-1: 0] frame_cube_flat
);

    always @(posedge clk) begin
        case(display_mode)
            `UART_MODE:     frame_cube_flat <= frame_valid_uart ? frame_cube_uart_flat : frame_cube_flat;
            `GEN_MODE:     frame_cube_flat <= frame_valid_default ? frame_cube_default_flat : frame_cube_flat;
            default:
                case(display_sel)
                    4'h0:   frame_cube_flat <= 256'hff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff;    //全亮
                    4'h1:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_ff_ff_ff_ff_ff_ff_ff_ff;    //1层
                    4'h2:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_ff_ff_ff_ff_ff_ff_ff_ff_00_00_00_00_00_00_00_00;    //2
                    4'h3:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_ff_ff_ff_ff_ff_ff_ff_ff_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;    //3
                    4'h4:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_ff_ff_ff_ff_ff_ff_ff_ff_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;    //4
                    4'h5:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_ff_ff_ff_ff_ff_ff_ff_ff_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;    //5
                    4'h6:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_ff_ff_ff_ff_ff_ff_ff_ff_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;    //6
                    4'h7:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_ff_ff_ff_ff_ff_ff_ff_ff_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;    //7
                    4'h8:   frame_cube_flat <= 256'hff_ff_ff_ff_ff_ff_ff_ff_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;    //8
                    4'h9:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_ff;    //1列
                    4'ha:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_ff_00;    //2
                    4'hb:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_ff_00_00;    //3
                    4'hc:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_01_01_01_01_01_01_01_01;    //1行
                    4'hd:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_01_01_01_01_01_01_01_01_00_00_00_00_00_00_00_00;    //2
                    4'he:   frame_cube_flat <= 256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_01_01_01_01_01_01_01_01_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00;    //3

                    4'hf:   frame_cube_flat <= 256'hff_81_81_81_81_81_81_ff_81_00_00_00_00_00_00_81_81_00_00_00_00_00_00_81_81_00_00_00_00_00_00_81_81_00_00_00_00_00_00_81_81_00_00_00_00_00_00_81_81_00_00_00_00_00_00_81_ff_81_81_81_81_81_81_ff;    //边框
                    // default: frame_cube_flat <= 256'hff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff_ff;
                endcase
        endcase
    end

    always @(posedge clk) begin
        if(rst) begin
            frame_cnt <= 0;
        end
        else if(frame_valid_uart | frame_valid_default)begin
            frame_cnt <= frame_cnt + 1;
        end
    end

endmodule