module uart_reciver (
    input wire clk,
    input wire rst,

    input wire rx,
    output wire tx, //no use
    output reg [7:0] frame_cube [63:0]
);
    
    
endmodule